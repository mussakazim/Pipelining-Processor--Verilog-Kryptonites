`timescale 1ns / 1ps


module AluMUX1(
    output [31:0] Mux1Output,
    input [31:0] RsData1
    );

     
	  assign Mux1Output = RsData1;

 
endmodule
